
module elc3_soc (
	clk_clk,
	reset_reset_n,
	sdram_clk_clk);	

	input		clk_clk;
	input		reset_reset_n;
	output		sdram_clk_clk;
endmodule
